package alu_pkg;

//standard UVM import & include

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "alu_transaction.sv"
`include "alu_config.sv"
`include "alu_sequence.sv"
`include "my_subscriber.sv"

endpackage: alu_pkg
